module identifica_cores 
(
    input wire       clock,
    input wire       reset,
    input wire       iniciar,
    input wire       pixel,
    output wire      addr_linha,
    output wire      addr_coluna,
    output wire      we,
    output wire [2:0] cor
);

endmodule